magic
tech sky130A
magscale 1 2
timestamp 1740732004
<< metal2 >>
rect 6510 8646 6566 9124
rect 6814 8642 6870 9108
rect 7118 8630 7174 9104
rect 7962 8828 8018 9124
rect 7858 8772 8018 8828
rect 7858 8616 7914 8772
rect 8346 8686 8402 9120
rect 8730 8690 8786 9116
rect 9294 8690 9350 9102
rect 8288 8630 8402 8686
rect 8680 8634 8786 8690
rect 9226 8634 9350 8690
rect 9598 8628 9654 9124
rect 9902 8684 9958 9116
rect 9834 8628 9958 8684
rect 10946 8694 11002 9124
rect 10946 8638 11062 8694
rect 11130 8638 11186 9104
rect 11314 8646 11370 9110
rect 11498 8638 11554 9110
rect 11682 8640 11738 9100
rect 11866 8696 11922 9098
rect 11816 8640 11922 8696
rect 16170 8646 16226 9124
rect 16474 8642 16530 9108
rect 16778 8630 16834 9104
rect 17622 8828 17678 9124
rect 17518 8772 17678 8828
rect 17518 8616 17574 8772
rect 18006 8686 18062 9120
rect 18390 8690 18446 9116
rect 18954 8690 19010 9102
rect 17948 8630 18062 8686
rect 18340 8634 18446 8690
rect 18886 8634 19010 8690
rect 19258 8628 19314 9124
rect 19562 8684 19618 9116
rect 19494 8628 19618 8684
rect 20606 8694 20662 9124
rect 20606 8638 20722 8694
rect 20790 8638 20846 9104
rect 20974 8646 21030 9110
rect 21158 8638 21214 9110
rect 21342 8640 21398 9100
rect 21526 8696 21582 9098
rect 21476 8640 21582 8696
rect 25830 8646 25886 9124
rect 26134 8642 26190 9108
rect 26438 8630 26494 9104
rect 27282 8828 27338 9124
rect 27178 8772 27338 8828
rect 27178 8616 27234 8772
rect 27666 8686 27722 9120
rect 28050 8690 28106 9116
rect 28614 8690 28670 9102
rect 27608 8630 27722 8686
rect 28000 8634 28106 8690
rect 28546 8634 28670 8690
rect 28918 8628 28974 9124
rect 29222 8684 29278 9116
rect 29154 8628 29278 8684
rect 30266 8694 30322 9124
rect 30266 8638 30382 8694
rect 30450 8638 30506 9104
rect 30634 8646 30690 9110
rect 30818 8638 30874 9110
rect 31002 8640 31058 9100
rect 31186 8696 31242 9098
rect 31136 8640 31242 8696
<< metal3 >>
rect 1521 6654 1919 6659
rect 194 6254 200 6654
rect 600 6653 1920 6654
rect 600 6255 1521 6653
rect 1919 6255 1920 6653
rect 600 6254 1920 6255
rect 1521 6249 1919 6254
rect 21123 3299 21413 3305
rect 11427 2971 11433 3289
rect 11751 2971 11757 3289
rect 21123 3003 21413 3009
rect 30780 2964 30786 3240
rect 31062 2964 31068 3240
<< via3 >>
rect 200 6254 600 6654
rect 1521 6255 1919 6653
rect 11433 2971 11751 3289
rect 21123 3009 21413 3299
rect 30786 2964 31062 3240
<< metal4 >>
rect 6134 44952 6194 45152
rect 6686 44952 6746 45152
rect 7238 44952 7298 45152
rect 7790 44952 7850 45152
rect 8342 44952 8402 45152
rect 8894 44952 8954 45152
rect 9446 44952 9506 45152
rect 9998 44952 10058 45152
rect 10550 44952 10610 45152
rect 11102 44952 11162 45152
rect 11654 44952 11714 45152
rect 12206 44952 12266 45152
rect 12758 44952 12818 45152
rect 13310 44952 13370 45152
rect 13862 44952 13922 45152
rect 14414 44952 14474 45152
rect 14966 44952 15026 45152
rect 15518 44952 15578 45152
rect 16070 44952 16130 45152
rect 16622 44952 16682 45152
rect 17174 44952 17234 45152
rect 17726 44952 17786 45152
rect 18278 44952 18338 45152
rect 18830 44952 18890 45152
rect 19382 44952 19442 45152
rect 19934 44952 19994 45152
rect 20486 44952 20546 45152
rect 21038 44952 21098 45152
rect 21590 44952 21650 45152
rect 22142 44952 22202 45152
rect 22694 44952 22754 45152
rect 23246 44952 23306 45152
rect 23798 44952 23858 45152
rect 24350 44952 24410 45152
rect 24902 44952 24962 45152
rect 25454 44952 25514 45152
rect 26006 44952 26066 45152
rect 26558 44952 26618 45152
rect 27110 44952 27170 45152
rect 27662 44952 27722 45152
rect 28214 44952 28274 45152
rect 28766 44952 28826 45152
rect 29318 44952 29378 45152
rect 200 6655 600 44152
rect 199 6654 601 6655
rect 199 6254 200 6654
rect 600 6254 601 6654
rect 199 6253 601 6254
rect 200 1000 600 6253
rect 800 6134 1200 44152
rect 1520 6653 25558 6654
rect 1520 6255 1521 6653
rect 1919 6255 25558 6653
rect 1520 6254 25558 6255
rect 800 5734 25558 6134
rect 800 1000 1200 5734
rect 21122 3299 24120 3300
rect 11432 3289 11752 3290
rect 11432 2971 11433 3289
rect 11751 2971 11752 3289
rect 21122 3009 21123 3299
rect 21413 3009 24120 3299
rect 21122 3008 24120 3009
rect 30785 3240 31063 3241
rect 11432 1916 11752 2971
rect 23884 2218 24064 3008
rect 30785 2964 30786 3240
rect 31062 2964 31063 3240
rect 23884 2038 26678 2218
rect 11432 1736 22814 1916
rect 11432 1666 11752 1736
rect 3314 0 3494 200
rect 7178 0 7358 200
rect 11042 0 11222 200
rect 14906 0 15086 200
rect 18770 0 18950 200
rect 22634 0 22814 1736
rect 26498 0 26678 2038
rect 30785 1634 31063 2964
rect 30362 1454 31063 1634
rect 30362 0 30542 1454
rect 30785 1405 31063 1454
rect 65000 1000 65400 44152
rect 65600 1000 66000 44152
use analog_control_wrapper  analog_control_wrapper_1
timestamp 1740731205
transform 1 0 2072 0 1 2042
box 514 496 62414 41000
use segdac  segdac_0
timestamp 1725599052
transform 1 0 27099 0 1 3114
box -1901 -360 4160 5600
use segdac  segdac_blue
timestamp 1725599052
transform 1 0 7779 0 1 3114
box -1901 -360 4160 5600
use segdac  segdac_green
timestamp 1725599052
transform 1 0 17439 0 1 3114
box -1901 -360 4160 5600
<< labels >>
flabel metal4 s 28766 44952 28826 45152 0 FreeSans 480 90 0 0 clk
port 0 nsew signal input
flabel metal4 s 29318 44952 29378 45152 0 FreeSans 480 90 0 0 ena
port 1 nsew signal input
flabel metal4 s 28214 44952 28274 45152 0 FreeSans 480 90 0 0 rst_n
port 2 nsew signal input
flabel metal4 s 30362 0 30542 200 0 FreeSans 960 0 0 0 ua[0]
port 3 nsew signal bidirectional
flabel metal4 s 26498 0 26678 200 0 FreeSans 960 0 0 0 ua[1]
port 4 nsew signal bidirectional
flabel metal4 s 22634 0 22814 200 0 FreeSans 960 0 0 0 ua[2]
port 5 nsew signal bidirectional
flabel metal4 s 18770 0 18950 200 0 FreeSans 960 0 0 0 ua[3]
port 6 nsew signal bidirectional
flabel metal4 s 14906 0 15086 200 0 FreeSans 960 0 0 0 ua[4]
port 7 nsew signal bidirectional
flabel metal4 s 11042 0 11222 200 0 FreeSans 960 0 0 0 ua[5]
port 8 nsew signal bidirectional
flabel metal4 s 7178 0 7358 200 0 FreeSans 960 0 0 0 ua[6]
port 9 nsew signal bidirectional
flabel metal4 s 3314 0 3494 200 0 FreeSans 960 0 0 0 ua[7]
port 10 nsew signal bidirectional
flabel metal4 s 27662 44952 27722 45152 0 FreeSans 480 90 0 0 ui_in[0]
port 11 nsew signal input
flabel metal4 s 27110 44952 27170 45152 0 FreeSans 480 90 0 0 ui_in[1]
port 12 nsew signal input
flabel metal4 s 26558 44952 26618 45152 0 FreeSans 480 90 0 0 ui_in[2]
port 13 nsew signal input
flabel metal4 s 26006 44952 26066 45152 0 FreeSans 480 90 0 0 ui_in[3]
port 14 nsew signal input
flabel metal4 s 25454 44952 25514 45152 0 FreeSans 480 90 0 0 ui_in[4]
port 15 nsew signal input
flabel metal4 s 24902 44952 24962 45152 0 FreeSans 480 90 0 0 ui_in[5]
port 16 nsew signal input
flabel metal4 s 24350 44952 24410 45152 0 FreeSans 480 90 0 0 ui_in[6]
port 17 nsew signal input
flabel metal4 s 23798 44952 23858 45152 0 FreeSans 480 90 0 0 ui_in[7]
port 18 nsew signal input
flabel metal4 s 23246 44952 23306 45152 0 FreeSans 480 90 0 0 uio_in[0]
port 19 nsew signal input
flabel metal4 s 22694 44952 22754 45152 0 FreeSans 480 90 0 0 uio_in[1]
port 20 nsew signal input
flabel metal4 s 22142 44952 22202 45152 0 FreeSans 480 90 0 0 uio_in[2]
port 21 nsew signal input
flabel metal4 s 21590 44952 21650 45152 0 FreeSans 480 90 0 0 uio_in[3]
port 22 nsew signal input
flabel metal4 s 21038 44952 21098 45152 0 FreeSans 480 90 0 0 uio_in[4]
port 23 nsew signal input
flabel metal4 s 20486 44952 20546 45152 0 FreeSans 480 90 0 0 uio_in[5]
port 24 nsew signal input
flabel metal4 s 19934 44952 19994 45152 0 FreeSans 480 90 0 0 uio_in[6]
port 25 nsew signal input
flabel metal4 s 19382 44952 19442 45152 0 FreeSans 480 90 0 0 uio_in[7]
port 26 nsew signal input
flabel metal4 s 9998 44952 10058 45152 0 FreeSans 480 90 0 0 uio_oe[0]
port 27 nsew signal output
flabel metal4 s 9446 44952 9506 45152 0 FreeSans 480 90 0 0 uio_oe[1]
port 28 nsew signal output
flabel metal4 s 8894 44952 8954 45152 0 FreeSans 480 90 0 0 uio_oe[2]
port 29 nsew signal output
flabel metal4 s 8342 44952 8402 45152 0 FreeSans 480 90 0 0 uio_oe[3]
port 30 nsew signal output
flabel metal4 s 7790 44952 7850 45152 0 FreeSans 480 90 0 0 uio_oe[4]
port 31 nsew signal output
flabel metal4 s 7238 44952 7298 45152 0 FreeSans 480 90 0 0 uio_oe[5]
port 32 nsew signal output
flabel metal4 s 6686 44952 6746 45152 0 FreeSans 480 90 0 0 uio_oe[6]
port 33 nsew signal output
flabel metal4 s 6134 44952 6194 45152 0 FreeSans 480 90 0 0 uio_oe[7]
port 34 nsew signal output
flabel metal4 s 14414 44952 14474 45152 0 FreeSans 480 90 0 0 uio_out[0]
port 35 nsew signal output
flabel metal4 s 13862 44952 13922 45152 0 FreeSans 480 90 0 0 uio_out[1]
port 36 nsew signal output
flabel metal4 s 13310 44952 13370 45152 0 FreeSans 480 90 0 0 uio_out[2]
port 37 nsew signal output
flabel metal4 s 12758 44952 12818 45152 0 FreeSans 480 90 0 0 uio_out[3]
port 38 nsew signal output
flabel metal4 s 12206 44952 12266 45152 0 FreeSans 480 90 0 0 uio_out[4]
port 39 nsew signal output
flabel metal4 s 11654 44952 11714 45152 0 FreeSans 480 90 0 0 uio_out[5]
port 40 nsew signal output
flabel metal4 s 11102 44952 11162 45152 0 FreeSans 480 90 0 0 uio_out[6]
port 41 nsew signal output
flabel metal4 s 10550 44952 10610 45152 0 FreeSans 480 90 0 0 uio_out[7]
port 42 nsew signal output
flabel metal4 s 18830 44952 18890 45152 0 FreeSans 480 90 0 0 uo_out[0]
port 43 nsew signal output
flabel metal4 s 18278 44952 18338 45152 0 FreeSans 480 90 0 0 uo_out[1]
port 44 nsew signal output
flabel metal4 s 17726 44952 17786 45152 0 FreeSans 480 90 0 0 uo_out[2]
port 45 nsew signal output
flabel metal4 s 17174 44952 17234 45152 0 FreeSans 480 90 0 0 uo_out[3]
port 46 nsew signal output
flabel metal4 s 16622 44952 16682 45152 0 FreeSans 480 90 0 0 uo_out[4]
port 47 nsew signal output
flabel metal4 s 16070 44952 16130 45152 0 FreeSans 480 90 0 0 uo_out[5]
port 48 nsew signal output
flabel metal4 s 15518 44952 15578 45152 0 FreeSans 480 90 0 0 uo_out[6]
port 49 nsew signal output
flabel metal4 s 14966 44952 15026 45152 0 FreeSans 480 90 0 0 uo_out[7]
port 50 nsew signal output
flabel metal4 200 1000 600 44152 1 FreeSans 400 0 0 0 VDPWR
port 51 nsew power bidirectional
flabel metal4 800 1000 1200 44152 1 FreeSans 400 0 0 0 VGND
port 52 nsew ground bidirectional
flabel metal4 65000 1000 65400 44152 1 FreeSans 400 0 0 0 VDPWR
port 51 nsew power bidirectional
flabel metal4 65600 1000 66000 44152 1 FreeSans 400 0 0 0 VGND
port 52 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 66976 45152
<< end >>
