magic
tech sky130A
magscale 1 2
timestamp 1740794342
<< metal1 >>
rect 5810 5410 6090 5590
rect 5810 5120 5990 5410
rect 5780 5090 6020 5120
rect 5780 4910 5810 5090
rect 5990 4910 6020 5090
rect 5780 4880 6020 4910
<< via1 >>
rect 5810 4910 5990 5090
<< metal2 >>
rect 6120 44784 6210 44800
rect 6120 44728 6136 44784
rect 6192 44728 6210 44784
rect 6120 44710 6210 44728
rect 6672 44784 6762 44800
rect 6672 44728 6688 44784
rect 6744 44728 6762 44784
rect 6672 44710 6762 44728
rect 7224 44784 7314 44800
rect 7224 44728 7240 44784
rect 7296 44728 7314 44784
rect 7224 44710 7314 44728
rect 7776 44784 7866 44800
rect 7776 44728 7792 44784
rect 7848 44728 7866 44784
rect 7776 44710 7866 44728
rect 8328 44784 8418 44800
rect 8328 44728 8344 44784
rect 8400 44728 8418 44784
rect 8328 44710 8418 44728
rect 8880 44784 8970 44800
rect 8880 44728 8896 44784
rect 8952 44728 8970 44784
rect 8880 44710 8970 44728
rect 9432 44784 9522 44800
rect 9432 44728 9448 44784
rect 9504 44728 9522 44784
rect 9432 44710 9522 44728
rect 9984 44784 10074 44800
rect 9984 44728 10000 44784
rect 10056 44728 10074 44784
rect 9984 44710 10074 44728
rect 10536 44784 10626 44800
rect 10536 44728 10552 44784
rect 10608 44728 10626 44784
rect 10536 44710 10626 44728
rect 11088 44784 11178 44800
rect 11088 44728 11104 44784
rect 11160 44728 11178 44784
rect 11088 44710 11178 44728
rect 11640 44784 11730 44800
rect 11640 44728 11656 44784
rect 11712 44728 11730 44784
rect 11640 44710 11730 44728
rect 12192 44784 12282 44800
rect 12192 44728 12208 44784
rect 12264 44728 12282 44784
rect 12192 44710 12282 44728
rect 12744 44784 12834 44800
rect 12744 44728 12760 44784
rect 12816 44728 12834 44784
rect 12744 44710 12834 44728
rect 13296 44784 13386 44800
rect 13296 44728 13312 44784
rect 13368 44728 13386 44784
rect 13296 44710 13386 44728
rect 13848 44784 13938 44800
rect 13848 44728 13864 44784
rect 13920 44728 13938 44784
rect 13848 44710 13938 44728
rect 14400 44784 14490 44800
rect 14400 44728 14416 44784
rect 14472 44728 14490 44784
rect 14400 44710 14490 44728
rect 14952 44784 15042 44800
rect 14952 44728 14968 44784
rect 15024 44728 15042 44784
rect 14952 44710 15042 44728
rect 15504 44784 15594 44800
rect 15504 44728 15520 44784
rect 15576 44728 15594 44784
rect 15504 44710 15594 44728
rect 16056 44784 16146 44800
rect 16056 44728 16072 44784
rect 16128 44728 16146 44784
rect 16056 44710 16146 44728
rect 16608 44784 16698 44800
rect 16608 44728 16624 44784
rect 16680 44728 16698 44784
rect 16608 44710 16698 44728
rect 17160 44784 17250 44800
rect 17160 44728 17176 44784
rect 17232 44728 17250 44784
rect 17160 44710 17250 44728
rect 17712 44784 17802 44800
rect 17712 44728 17728 44784
rect 17784 44728 17802 44784
rect 17712 44710 17802 44728
rect 18264 44784 18354 44800
rect 18264 44728 18280 44784
rect 18336 44728 18354 44784
rect 18264 44710 18354 44728
rect 18816 44784 18906 44800
rect 18816 44728 18832 44784
rect 18888 44728 18906 44784
rect 18816 44710 18906 44728
rect 19368 44784 19458 44800
rect 19368 44728 19384 44784
rect 19440 44728 19458 44784
rect 19368 44710 19458 44728
rect 19920 44784 20010 44800
rect 19920 44728 19936 44784
rect 19992 44728 20010 44784
rect 19920 44710 20010 44728
rect 20472 44784 20562 44800
rect 20472 44728 20488 44784
rect 20544 44728 20562 44784
rect 20472 44710 20562 44728
rect 21024 44784 21114 44800
rect 21024 44728 21040 44784
rect 21096 44728 21114 44784
rect 21024 44710 21114 44728
rect 21576 44784 21666 44800
rect 21576 44728 21592 44784
rect 21648 44728 21666 44784
rect 21576 44710 21666 44728
rect 22128 44784 22218 44800
rect 22128 44728 22144 44784
rect 22200 44728 22218 44784
rect 22128 44710 22218 44728
rect 22680 44784 22770 44800
rect 22680 44728 22696 44784
rect 22752 44728 22770 44784
rect 22680 44710 22770 44728
rect 23232 44784 23322 44800
rect 23232 44728 23248 44784
rect 23304 44728 23322 44784
rect 23232 44710 23322 44728
rect 23784 44784 23874 44800
rect 23784 44728 23800 44784
rect 23856 44728 23874 44784
rect 23784 44710 23874 44728
rect 24336 44784 24426 44800
rect 24336 44728 24352 44784
rect 24408 44728 24426 44784
rect 24336 44710 24426 44728
rect 24888 44784 24978 44800
rect 24888 44728 24904 44784
rect 24960 44728 24978 44784
rect 24888 44710 24978 44728
rect 25440 44784 25530 44800
rect 25440 44728 25456 44784
rect 25512 44728 25530 44784
rect 25440 44710 25530 44728
rect 25992 44784 26082 44800
rect 25992 44728 26008 44784
rect 26064 44728 26082 44784
rect 25992 44710 26082 44728
rect 26544 44784 26634 44800
rect 26544 44728 26560 44784
rect 26616 44728 26634 44784
rect 26544 44710 26634 44728
rect 27096 44784 27186 44800
rect 27096 44728 27112 44784
rect 27168 44728 27186 44784
rect 27096 44710 27186 44728
rect 27648 44784 27738 44800
rect 27648 44728 27664 44784
rect 27720 44728 27738 44784
rect 27648 44710 27738 44728
rect 28200 44784 28290 44800
rect 28200 44728 28216 44784
rect 28272 44728 28290 44784
rect 28200 44710 28290 44728
rect 28752 44784 28842 44800
rect 28752 44728 28768 44784
rect 28824 44728 28842 44784
rect 28752 44710 28842 44728
rect 29304 44784 29394 44800
rect 29304 44728 29320 44784
rect 29376 44728 29394 44784
rect 29304 44710 29394 44728
rect 6134 44532 6194 44710
rect 6686 44532 6746 44710
rect 7238 44532 7298 44710
rect 7790 44532 7850 44710
rect 8342 44532 8402 44710
rect 8894 44532 8954 44710
rect 9446 44532 9506 44710
rect 9998 44532 10058 44710
rect 10550 44532 10610 44710
rect 11102 44532 11162 44710
rect 11654 44532 11714 44710
rect 12206 44532 12266 44710
rect 12758 44532 12818 44710
rect 13310 44532 13370 44710
rect 13862 44532 13922 44710
rect 14414 44532 14474 44710
rect 14966 44532 15026 44710
rect 15518 44532 15578 44710
rect 16070 44532 16130 44710
rect 16622 44532 16682 44710
rect 17174 44532 17234 44710
rect 17726 44532 17786 44710
rect 18278 44532 18338 44710
rect 18830 44532 18890 44710
rect 19382 44532 19442 44710
rect 19934 44532 19994 44710
rect 20486 44532 20546 44710
rect 21038 44532 21098 44710
rect 21590 44532 21650 44710
rect 22142 44532 22202 44710
rect 22694 44532 22754 44710
rect 23246 44532 23306 44710
rect 23798 44532 23858 44710
rect 24350 44532 24410 44710
rect 24902 44532 24962 44710
rect 25454 44532 25514 44710
rect 26006 44532 26066 44710
rect 26558 44532 26618 44710
rect 27110 44532 27170 44710
rect 27662 44532 27722 44710
rect 28214 44532 28274 44710
rect 28766 44532 28826 44710
rect 29318 44532 29378 44710
rect 6138 42996 6194 44532
rect 6690 42996 6746 44532
rect 7242 42996 7298 44532
rect 7794 42996 7850 44532
rect 8346 42996 8402 44532
rect 8898 42996 8954 44532
rect 9450 42996 9506 44532
rect 10002 42996 10058 44532
rect 10554 42996 10610 44532
rect 11106 42996 11162 44532
rect 11658 42996 11714 44532
rect 12210 42996 12266 44532
rect 12762 42996 12818 44532
rect 13314 42996 13370 44532
rect 13866 42996 13922 44532
rect 14418 42996 14474 44532
rect 14970 42996 15026 44532
rect 15522 42996 15578 44532
rect 16074 42996 16130 44532
rect 16626 42996 16682 44532
rect 17178 42996 17234 44532
rect 17730 42996 17786 44532
rect 18282 42996 18338 44532
rect 18834 42996 18890 44532
rect 19386 42996 19442 44532
rect 19938 42996 19994 44532
rect 20490 42996 20546 44532
rect 21042 42996 21098 44532
rect 21594 42996 21650 44532
rect 22146 42996 22202 44532
rect 22698 42996 22754 44532
rect 23250 42996 23306 44532
rect 23802 42996 23858 44532
rect 24354 42996 24410 44532
rect 24906 42996 24962 44532
rect 25458 42996 25514 44532
rect 26010 42996 26066 44532
rect 26562 42996 26618 44532
rect 27114 42996 27170 44532
rect 27666 42996 27722 44532
rect 28218 42996 28274 44532
rect 28770 42996 28826 44532
rect 29322 42996 29378 44532
rect 6510 8646 6566 9124
rect 6814 8642 6870 9108
rect 7118 8630 7174 9104
rect 7962 8828 8018 9124
rect 7858 8772 8018 8828
rect 7858 8616 7914 8772
rect 8346 8686 8402 9120
rect 8730 8690 8786 9116
rect 9294 8690 9350 9102
rect 8288 8630 8402 8686
rect 8680 8634 8786 8690
rect 9226 8634 9350 8690
rect 9598 8628 9654 9124
rect 9902 8684 9958 9116
rect 9834 8628 9958 8684
rect 10946 8694 11002 9124
rect 10946 8638 11062 8694
rect 11130 8638 11186 9104
rect 11314 8646 11370 9110
rect 11498 8638 11554 9110
rect 11682 8640 11738 9100
rect 11866 8696 11922 9098
rect 11816 8640 11922 8696
rect 16170 8646 16226 9124
rect 16474 8642 16530 9108
rect 16778 8630 16834 9104
rect 17622 8828 17678 9124
rect 17518 8772 17678 8828
rect 17518 8616 17574 8772
rect 18006 8686 18062 9120
rect 18390 8690 18446 9116
rect 18954 8690 19010 9102
rect 17948 8630 18062 8686
rect 18340 8634 18446 8690
rect 18886 8634 19010 8690
rect 19258 8628 19314 9124
rect 19562 8684 19618 9116
rect 19494 8628 19618 8684
rect 20606 8694 20662 9124
rect 20606 8638 20722 8694
rect 20790 8638 20846 9104
rect 20974 8646 21030 9110
rect 21158 8638 21214 9110
rect 21342 8640 21398 9100
rect 21526 8696 21582 9098
rect 21476 8640 21582 8696
rect 25830 8646 25886 9124
rect 26134 8642 26190 9108
rect 26438 8630 26494 9104
rect 27282 8828 27338 9124
rect 27178 8772 27338 8828
rect 27178 8616 27234 8772
rect 27666 8686 27722 9120
rect 28050 8690 28106 9116
rect 28614 8690 28670 9102
rect 27608 8630 27722 8686
rect 28000 8634 28106 8690
rect 28546 8634 28670 8690
rect 28918 8628 28974 9124
rect 29222 8684 29278 9116
rect 29154 8628 29278 8684
rect 30266 8694 30322 9124
rect 30266 8638 30382 8694
rect 30450 8638 30506 9104
rect 30634 8646 30690 9110
rect 30818 8638 30874 9110
rect 31002 8640 31058 9100
rect 31186 8696 31242 9098
rect 31136 8640 31242 8696
rect 5780 5090 6020 5120
rect 5780 4910 5810 5090
rect 5990 4910 6020 5090
rect 5780 4880 6020 4910
<< via2 >>
rect 6136 44728 6192 44784
rect 6688 44728 6744 44784
rect 7240 44728 7296 44784
rect 7792 44728 7848 44784
rect 8344 44728 8400 44784
rect 8896 44728 8952 44784
rect 9448 44728 9504 44784
rect 10000 44728 10056 44784
rect 10552 44728 10608 44784
rect 11104 44728 11160 44784
rect 11656 44728 11712 44784
rect 12208 44728 12264 44784
rect 12760 44728 12816 44784
rect 13312 44728 13368 44784
rect 13864 44728 13920 44784
rect 14416 44728 14472 44784
rect 14968 44728 15024 44784
rect 15520 44728 15576 44784
rect 16072 44728 16128 44784
rect 16624 44728 16680 44784
rect 17176 44728 17232 44784
rect 17728 44728 17784 44784
rect 18280 44728 18336 44784
rect 18832 44728 18888 44784
rect 19384 44728 19440 44784
rect 19936 44728 19992 44784
rect 20488 44728 20544 44784
rect 21040 44728 21096 44784
rect 21592 44728 21648 44784
rect 22144 44728 22200 44784
rect 22696 44728 22752 44784
rect 23248 44728 23304 44784
rect 23800 44728 23856 44784
rect 24352 44728 24408 44784
rect 24904 44728 24960 44784
rect 25456 44728 25512 44784
rect 26008 44728 26064 44784
rect 26560 44728 26616 44784
rect 27112 44728 27168 44784
rect 27664 44728 27720 44784
rect 28216 44728 28272 44784
rect 28768 44728 28824 44784
rect 29320 44728 29376 44784
rect 5815 4915 5985 5085
<< metal3 >>
rect 6110 44788 6220 44810
rect 6110 44724 6132 44788
rect 6196 44724 6220 44788
rect 6110 44700 6220 44724
rect 6662 44788 6772 44810
rect 6662 44724 6684 44788
rect 6748 44724 6772 44788
rect 6662 44700 6772 44724
rect 7214 44788 7324 44810
rect 7214 44724 7236 44788
rect 7300 44724 7324 44788
rect 7214 44700 7324 44724
rect 7766 44788 7876 44810
rect 7766 44724 7788 44788
rect 7852 44724 7876 44788
rect 7766 44700 7876 44724
rect 8318 44788 8428 44810
rect 8318 44724 8340 44788
rect 8404 44724 8428 44788
rect 8318 44700 8428 44724
rect 8870 44788 8980 44810
rect 8870 44724 8892 44788
rect 8956 44724 8980 44788
rect 8870 44700 8980 44724
rect 9422 44788 9532 44810
rect 9422 44724 9444 44788
rect 9508 44724 9532 44788
rect 9422 44700 9532 44724
rect 9974 44788 10084 44810
rect 9974 44724 9996 44788
rect 10060 44724 10084 44788
rect 9974 44700 10084 44724
rect 10526 44788 10636 44810
rect 10526 44724 10548 44788
rect 10612 44724 10636 44788
rect 10526 44700 10636 44724
rect 11078 44788 11188 44810
rect 11078 44724 11100 44788
rect 11164 44724 11188 44788
rect 11078 44700 11188 44724
rect 11630 44788 11740 44810
rect 11630 44724 11652 44788
rect 11716 44724 11740 44788
rect 11630 44700 11740 44724
rect 12182 44788 12292 44810
rect 12182 44724 12204 44788
rect 12268 44724 12292 44788
rect 12182 44700 12292 44724
rect 12734 44788 12844 44810
rect 12734 44724 12756 44788
rect 12820 44724 12844 44788
rect 12734 44700 12844 44724
rect 13286 44788 13396 44810
rect 13286 44724 13308 44788
rect 13372 44724 13396 44788
rect 13286 44700 13396 44724
rect 13838 44788 13948 44810
rect 13838 44724 13860 44788
rect 13924 44724 13948 44788
rect 13838 44700 13948 44724
rect 14390 44788 14500 44810
rect 14390 44724 14412 44788
rect 14476 44724 14500 44788
rect 14390 44700 14500 44724
rect 14942 44788 15052 44810
rect 14942 44724 14964 44788
rect 15028 44724 15052 44788
rect 14942 44700 15052 44724
rect 15494 44788 15604 44810
rect 15494 44724 15516 44788
rect 15580 44724 15604 44788
rect 15494 44700 15604 44724
rect 16046 44788 16156 44810
rect 16046 44724 16068 44788
rect 16132 44724 16156 44788
rect 16046 44700 16156 44724
rect 16598 44788 16708 44810
rect 16598 44724 16620 44788
rect 16684 44724 16708 44788
rect 16598 44700 16708 44724
rect 17150 44788 17260 44810
rect 17150 44724 17172 44788
rect 17236 44724 17260 44788
rect 17150 44700 17260 44724
rect 17702 44788 17812 44810
rect 17702 44724 17724 44788
rect 17788 44724 17812 44788
rect 17702 44700 17812 44724
rect 18254 44788 18364 44810
rect 18254 44724 18276 44788
rect 18340 44724 18364 44788
rect 18254 44700 18364 44724
rect 18806 44788 18916 44810
rect 18806 44724 18828 44788
rect 18892 44724 18916 44788
rect 18806 44700 18916 44724
rect 19358 44788 19468 44810
rect 19358 44724 19380 44788
rect 19444 44724 19468 44788
rect 19358 44700 19468 44724
rect 19910 44788 20020 44810
rect 19910 44724 19932 44788
rect 19996 44724 20020 44788
rect 19910 44700 20020 44724
rect 20462 44788 20572 44810
rect 20462 44724 20484 44788
rect 20548 44724 20572 44788
rect 20462 44700 20572 44724
rect 21014 44788 21124 44810
rect 21014 44724 21036 44788
rect 21100 44724 21124 44788
rect 21014 44700 21124 44724
rect 21566 44788 21676 44810
rect 21566 44724 21588 44788
rect 21652 44724 21676 44788
rect 21566 44700 21676 44724
rect 22118 44788 22228 44810
rect 22118 44724 22140 44788
rect 22204 44724 22228 44788
rect 22118 44700 22228 44724
rect 22670 44788 22780 44810
rect 22670 44724 22692 44788
rect 22756 44724 22780 44788
rect 22670 44700 22780 44724
rect 23222 44788 23332 44810
rect 23222 44724 23244 44788
rect 23308 44724 23332 44788
rect 23222 44700 23332 44724
rect 23774 44788 23884 44810
rect 23774 44724 23796 44788
rect 23860 44724 23884 44788
rect 23774 44700 23884 44724
rect 24326 44788 24436 44810
rect 24326 44724 24348 44788
rect 24412 44724 24436 44788
rect 24326 44700 24436 44724
rect 24878 44788 24988 44810
rect 24878 44724 24900 44788
rect 24964 44724 24988 44788
rect 24878 44700 24988 44724
rect 25430 44788 25540 44810
rect 25430 44724 25452 44788
rect 25516 44724 25540 44788
rect 25430 44700 25540 44724
rect 25982 44788 26092 44810
rect 25982 44724 26004 44788
rect 26068 44724 26092 44788
rect 25982 44700 26092 44724
rect 26534 44788 26644 44810
rect 26534 44724 26556 44788
rect 26620 44724 26644 44788
rect 26534 44700 26644 44724
rect 27086 44788 27196 44810
rect 27086 44724 27108 44788
rect 27172 44724 27196 44788
rect 27086 44700 27196 44724
rect 27638 44788 27748 44810
rect 27638 44724 27660 44788
rect 27724 44724 27748 44788
rect 27638 44700 27748 44724
rect 28190 44788 28300 44810
rect 28190 44724 28212 44788
rect 28276 44724 28300 44788
rect 28190 44700 28300 44724
rect 28742 44788 28852 44810
rect 28742 44724 28764 44788
rect 28828 44724 28852 44788
rect 28742 44700 28852 44724
rect 29294 44788 29404 44810
rect 29294 44724 29316 44788
rect 29380 44724 29404 44788
rect 29294 44700 29404 44724
rect 4400 43300 5300 43400
rect 6300 43300 6800 43400
rect 14074 43300 14574 43400
rect 21848 43300 22348 43400
rect 29622 43300 30122 43400
rect 37396 43300 37896 43400
rect 45170 43300 45670 43400
rect 52944 43300 53444 43400
rect 60718 43300 61218 43400
rect 65600 43300 66100 43400
rect 4400 42800 4500 43300
rect 5200 42800 6400 43300
rect 6700 42800 14174 43300
rect 14474 42800 21948 43300
rect 22248 42800 29722 43300
rect 30022 42800 37496 43300
rect 37796 42800 45270 43300
rect 45570 42800 53044 43300
rect 53344 42800 60818 43300
rect 61118 42800 65700 43300
rect 66000 42800 66100 43300
rect 4400 42700 5300 42800
rect 6300 42700 6800 42800
rect 14074 42700 14574 42800
rect 21848 42700 22348 42800
rect 29622 42700 30122 42800
rect 37396 42700 37896 42800
rect 45170 42700 45670 42800
rect 52944 42700 53444 42800
rect 60718 42700 61218 42800
rect 65600 42700 66100 42800
rect 1521 6654 1919 6659
rect 194 6254 200 6654
rect 600 6653 1920 6654
rect 600 6255 1521 6653
rect 1919 6255 1920 6653
rect 600 6254 1920 6255
rect 1521 6249 1919 6254
rect 5780 5089 6020 5120
rect 5780 4911 5811 5089
rect 5989 4911 6020 5089
rect 5780 4880 6020 4911
rect 21123 3299 21413 3305
rect 11427 2971 11433 3289
rect 11751 2971 11757 3289
rect 21123 3003 21413 3009
rect 30780 2964 30786 3240
rect 31062 2964 31068 3240
<< via3 >>
rect 6132 44784 6196 44788
rect 6132 44728 6136 44784
rect 6136 44728 6192 44784
rect 6192 44728 6196 44784
rect 6132 44724 6196 44728
rect 6684 44784 6748 44788
rect 6684 44728 6688 44784
rect 6688 44728 6744 44784
rect 6744 44728 6748 44784
rect 6684 44724 6748 44728
rect 7236 44784 7300 44788
rect 7236 44728 7240 44784
rect 7240 44728 7296 44784
rect 7296 44728 7300 44784
rect 7236 44724 7300 44728
rect 7788 44784 7852 44788
rect 7788 44728 7792 44784
rect 7792 44728 7848 44784
rect 7848 44728 7852 44784
rect 7788 44724 7852 44728
rect 8340 44784 8404 44788
rect 8340 44728 8344 44784
rect 8344 44728 8400 44784
rect 8400 44728 8404 44784
rect 8340 44724 8404 44728
rect 8892 44784 8956 44788
rect 8892 44728 8896 44784
rect 8896 44728 8952 44784
rect 8952 44728 8956 44784
rect 8892 44724 8956 44728
rect 9444 44784 9508 44788
rect 9444 44728 9448 44784
rect 9448 44728 9504 44784
rect 9504 44728 9508 44784
rect 9444 44724 9508 44728
rect 9996 44784 10060 44788
rect 9996 44728 10000 44784
rect 10000 44728 10056 44784
rect 10056 44728 10060 44784
rect 9996 44724 10060 44728
rect 10548 44784 10612 44788
rect 10548 44728 10552 44784
rect 10552 44728 10608 44784
rect 10608 44728 10612 44784
rect 10548 44724 10612 44728
rect 11100 44784 11164 44788
rect 11100 44728 11104 44784
rect 11104 44728 11160 44784
rect 11160 44728 11164 44784
rect 11100 44724 11164 44728
rect 11652 44784 11716 44788
rect 11652 44728 11656 44784
rect 11656 44728 11712 44784
rect 11712 44728 11716 44784
rect 11652 44724 11716 44728
rect 12204 44784 12268 44788
rect 12204 44728 12208 44784
rect 12208 44728 12264 44784
rect 12264 44728 12268 44784
rect 12204 44724 12268 44728
rect 12756 44784 12820 44788
rect 12756 44728 12760 44784
rect 12760 44728 12816 44784
rect 12816 44728 12820 44784
rect 12756 44724 12820 44728
rect 13308 44784 13372 44788
rect 13308 44728 13312 44784
rect 13312 44728 13368 44784
rect 13368 44728 13372 44784
rect 13308 44724 13372 44728
rect 13860 44784 13924 44788
rect 13860 44728 13864 44784
rect 13864 44728 13920 44784
rect 13920 44728 13924 44784
rect 13860 44724 13924 44728
rect 14412 44784 14476 44788
rect 14412 44728 14416 44784
rect 14416 44728 14472 44784
rect 14472 44728 14476 44784
rect 14412 44724 14476 44728
rect 14964 44784 15028 44788
rect 14964 44728 14968 44784
rect 14968 44728 15024 44784
rect 15024 44728 15028 44784
rect 14964 44724 15028 44728
rect 15516 44784 15580 44788
rect 15516 44728 15520 44784
rect 15520 44728 15576 44784
rect 15576 44728 15580 44784
rect 15516 44724 15580 44728
rect 16068 44784 16132 44788
rect 16068 44728 16072 44784
rect 16072 44728 16128 44784
rect 16128 44728 16132 44784
rect 16068 44724 16132 44728
rect 16620 44784 16684 44788
rect 16620 44728 16624 44784
rect 16624 44728 16680 44784
rect 16680 44728 16684 44784
rect 16620 44724 16684 44728
rect 17172 44784 17236 44788
rect 17172 44728 17176 44784
rect 17176 44728 17232 44784
rect 17232 44728 17236 44784
rect 17172 44724 17236 44728
rect 17724 44784 17788 44788
rect 17724 44728 17728 44784
rect 17728 44728 17784 44784
rect 17784 44728 17788 44784
rect 17724 44724 17788 44728
rect 18276 44784 18340 44788
rect 18276 44728 18280 44784
rect 18280 44728 18336 44784
rect 18336 44728 18340 44784
rect 18276 44724 18340 44728
rect 18828 44784 18892 44788
rect 18828 44728 18832 44784
rect 18832 44728 18888 44784
rect 18888 44728 18892 44784
rect 18828 44724 18892 44728
rect 19380 44784 19444 44788
rect 19380 44728 19384 44784
rect 19384 44728 19440 44784
rect 19440 44728 19444 44784
rect 19380 44724 19444 44728
rect 19932 44784 19996 44788
rect 19932 44728 19936 44784
rect 19936 44728 19992 44784
rect 19992 44728 19996 44784
rect 19932 44724 19996 44728
rect 20484 44784 20548 44788
rect 20484 44728 20488 44784
rect 20488 44728 20544 44784
rect 20544 44728 20548 44784
rect 20484 44724 20548 44728
rect 21036 44784 21100 44788
rect 21036 44728 21040 44784
rect 21040 44728 21096 44784
rect 21096 44728 21100 44784
rect 21036 44724 21100 44728
rect 21588 44784 21652 44788
rect 21588 44728 21592 44784
rect 21592 44728 21648 44784
rect 21648 44728 21652 44784
rect 21588 44724 21652 44728
rect 22140 44784 22204 44788
rect 22140 44728 22144 44784
rect 22144 44728 22200 44784
rect 22200 44728 22204 44784
rect 22140 44724 22204 44728
rect 22692 44784 22756 44788
rect 22692 44728 22696 44784
rect 22696 44728 22752 44784
rect 22752 44728 22756 44784
rect 22692 44724 22756 44728
rect 23244 44784 23308 44788
rect 23244 44728 23248 44784
rect 23248 44728 23304 44784
rect 23304 44728 23308 44784
rect 23244 44724 23308 44728
rect 23796 44784 23860 44788
rect 23796 44728 23800 44784
rect 23800 44728 23856 44784
rect 23856 44728 23860 44784
rect 23796 44724 23860 44728
rect 24348 44784 24412 44788
rect 24348 44728 24352 44784
rect 24352 44728 24408 44784
rect 24408 44728 24412 44784
rect 24348 44724 24412 44728
rect 24900 44784 24964 44788
rect 24900 44728 24904 44784
rect 24904 44728 24960 44784
rect 24960 44728 24964 44784
rect 24900 44724 24964 44728
rect 25452 44784 25516 44788
rect 25452 44728 25456 44784
rect 25456 44728 25512 44784
rect 25512 44728 25516 44784
rect 25452 44724 25516 44728
rect 26004 44784 26068 44788
rect 26004 44728 26008 44784
rect 26008 44728 26064 44784
rect 26064 44728 26068 44784
rect 26004 44724 26068 44728
rect 26556 44784 26620 44788
rect 26556 44728 26560 44784
rect 26560 44728 26616 44784
rect 26616 44728 26620 44784
rect 26556 44724 26620 44728
rect 27108 44784 27172 44788
rect 27108 44728 27112 44784
rect 27112 44728 27168 44784
rect 27168 44728 27172 44784
rect 27108 44724 27172 44728
rect 27660 44784 27724 44788
rect 27660 44728 27664 44784
rect 27664 44728 27720 44784
rect 27720 44728 27724 44784
rect 27660 44724 27724 44728
rect 28212 44784 28276 44788
rect 28212 44728 28216 44784
rect 28216 44728 28272 44784
rect 28272 44728 28276 44784
rect 28212 44724 28276 44728
rect 28764 44784 28828 44788
rect 28764 44728 28768 44784
rect 28768 44728 28824 44784
rect 28824 44728 28828 44784
rect 28764 44724 28828 44728
rect 29316 44784 29380 44788
rect 29316 44728 29320 44784
rect 29320 44728 29376 44784
rect 29376 44728 29380 44784
rect 29316 44724 29380 44728
rect 4500 42800 5200 43300
rect 6400 42800 6700 43300
rect 14174 42800 14474 43300
rect 21948 42800 22248 43300
rect 29722 42800 30022 43300
rect 37496 42800 37796 43300
rect 45270 42800 45570 43300
rect 53044 42800 53344 43300
rect 60818 42800 61118 43300
rect 65700 42800 66000 43300
rect 200 6254 600 6654
rect 1521 6255 1919 6653
rect 5811 5085 5989 5089
rect 5811 4915 5815 5085
rect 5815 4915 5985 5085
rect 5985 4915 5989 5085
rect 5811 4911 5989 4915
rect 11433 2971 11751 3289
rect 21123 3009 21413 3299
rect 30786 2964 31062 3240
<< metal4 >>
rect 200 44400 2400 44900
rect 6134 44800 6194 45152
rect 6686 44800 6746 45152
rect 7238 44800 7298 45152
rect 7790 44800 7850 45152
rect 8342 44800 8402 45152
rect 8894 44800 8954 45152
rect 9446 44800 9506 45152
rect 9998 44800 10058 45152
rect 10550 44800 10610 45152
rect 11102 44800 11162 45152
rect 11654 44800 11714 45152
rect 12206 44800 12266 45152
rect 12758 44800 12818 45152
rect 13310 44800 13370 45152
rect 13862 44800 13922 45152
rect 14414 44800 14474 45152
rect 14966 44800 15026 45152
rect 15518 44800 15578 45152
rect 16070 44800 16130 45152
rect 16622 44800 16682 45152
rect 17174 44800 17234 45152
rect 17726 44800 17786 45152
rect 18278 44800 18338 45152
rect 18830 44800 18890 45152
rect 19382 44800 19442 45152
rect 19934 44800 19994 45152
rect 20486 44800 20546 45152
rect 21038 44800 21098 45152
rect 21590 44800 21650 45152
rect 22142 44800 22202 45152
rect 22694 44800 22754 45152
rect 23246 44800 23306 45152
rect 23798 44800 23858 45152
rect 24350 44800 24410 45152
rect 24902 44800 24962 45152
rect 25454 44800 25514 45152
rect 26006 44800 26066 45152
rect 26558 44800 26618 45152
rect 27110 44800 27170 45152
rect 27662 44800 27722 45152
rect 28214 44800 28274 45152
rect 28766 44800 28826 45152
rect 29318 44800 29378 45152
rect 6120 44788 6210 44800
rect 6120 44724 6132 44788
rect 6196 44724 6210 44788
rect 6120 44710 6210 44724
rect 6672 44788 6762 44800
rect 6672 44724 6684 44788
rect 6748 44724 6762 44788
rect 6672 44710 6762 44724
rect 7224 44788 7314 44800
rect 7224 44724 7236 44788
rect 7300 44724 7314 44788
rect 7224 44710 7314 44724
rect 7776 44788 7866 44800
rect 7776 44724 7788 44788
rect 7852 44724 7866 44788
rect 7776 44710 7866 44724
rect 8328 44788 8418 44800
rect 8328 44724 8340 44788
rect 8404 44724 8418 44788
rect 8328 44710 8418 44724
rect 8880 44788 8970 44800
rect 8880 44724 8892 44788
rect 8956 44724 8970 44788
rect 8880 44710 8970 44724
rect 9432 44788 9522 44800
rect 9432 44724 9444 44788
rect 9508 44724 9522 44788
rect 9432 44710 9522 44724
rect 9984 44788 10074 44800
rect 9984 44724 9996 44788
rect 10060 44724 10074 44788
rect 9984 44710 10074 44724
rect 10536 44788 10626 44800
rect 10536 44724 10548 44788
rect 10612 44724 10626 44788
rect 10536 44710 10626 44724
rect 11088 44788 11178 44800
rect 11088 44724 11100 44788
rect 11164 44724 11178 44788
rect 11088 44710 11178 44724
rect 11640 44788 11730 44800
rect 11640 44724 11652 44788
rect 11716 44724 11730 44788
rect 11640 44710 11730 44724
rect 12192 44788 12282 44800
rect 12192 44724 12204 44788
rect 12268 44724 12282 44788
rect 12192 44710 12282 44724
rect 12744 44788 12834 44800
rect 12744 44724 12756 44788
rect 12820 44724 12834 44788
rect 12744 44710 12834 44724
rect 13296 44788 13386 44800
rect 13296 44724 13308 44788
rect 13372 44724 13386 44788
rect 13296 44710 13386 44724
rect 13848 44788 13938 44800
rect 13848 44724 13860 44788
rect 13924 44724 13938 44788
rect 13848 44710 13938 44724
rect 14400 44788 14490 44800
rect 14400 44724 14412 44788
rect 14476 44724 14490 44788
rect 14400 44710 14490 44724
rect 14952 44788 15042 44800
rect 14952 44724 14964 44788
rect 15028 44724 15042 44788
rect 14952 44710 15042 44724
rect 15504 44788 15594 44800
rect 15504 44724 15516 44788
rect 15580 44724 15594 44788
rect 15504 44710 15594 44724
rect 16056 44788 16146 44800
rect 16056 44724 16068 44788
rect 16132 44724 16146 44788
rect 16056 44710 16146 44724
rect 16608 44788 16698 44800
rect 16608 44724 16620 44788
rect 16684 44724 16698 44788
rect 16608 44710 16698 44724
rect 17160 44788 17250 44800
rect 17160 44724 17172 44788
rect 17236 44724 17250 44788
rect 17160 44710 17250 44724
rect 17712 44788 17802 44800
rect 17712 44724 17724 44788
rect 17788 44724 17802 44788
rect 17712 44710 17802 44724
rect 18264 44788 18354 44800
rect 18264 44724 18276 44788
rect 18340 44724 18354 44788
rect 18264 44710 18354 44724
rect 18816 44788 18906 44800
rect 18816 44724 18828 44788
rect 18892 44724 18906 44788
rect 18816 44710 18906 44724
rect 19368 44788 19458 44800
rect 19368 44724 19380 44788
rect 19444 44724 19458 44788
rect 19368 44710 19458 44724
rect 19920 44788 20010 44800
rect 19920 44724 19932 44788
rect 19996 44724 20010 44788
rect 19920 44710 20010 44724
rect 20472 44788 20562 44800
rect 20472 44724 20484 44788
rect 20548 44724 20562 44788
rect 20472 44710 20562 44724
rect 21024 44788 21114 44800
rect 21024 44724 21036 44788
rect 21100 44724 21114 44788
rect 21024 44710 21114 44724
rect 21576 44788 21666 44800
rect 21576 44724 21588 44788
rect 21652 44724 21666 44788
rect 21576 44710 21666 44724
rect 22128 44788 22218 44800
rect 22128 44724 22140 44788
rect 22204 44724 22218 44788
rect 22128 44710 22218 44724
rect 22680 44788 22770 44800
rect 22680 44724 22692 44788
rect 22756 44724 22770 44788
rect 22680 44710 22770 44724
rect 23232 44788 23322 44800
rect 23232 44724 23244 44788
rect 23308 44724 23322 44788
rect 23232 44710 23322 44724
rect 23784 44788 23874 44800
rect 23784 44724 23796 44788
rect 23860 44724 23874 44788
rect 23784 44710 23874 44724
rect 24336 44788 24426 44800
rect 24336 44724 24348 44788
rect 24412 44724 24426 44788
rect 24336 44710 24426 44724
rect 24888 44788 24978 44800
rect 24888 44724 24900 44788
rect 24964 44724 24978 44788
rect 24888 44710 24978 44724
rect 25440 44788 25530 44800
rect 25440 44724 25452 44788
rect 25516 44724 25530 44788
rect 25440 44710 25530 44724
rect 25992 44788 26082 44800
rect 25992 44724 26004 44788
rect 26068 44724 26082 44788
rect 25992 44710 26082 44724
rect 26544 44788 26634 44800
rect 26544 44724 26556 44788
rect 26620 44724 26634 44788
rect 26544 44710 26634 44724
rect 27096 44788 27186 44800
rect 27096 44724 27108 44788
rect 27172 44724 27186 44788
rect 27096 44710 27186 44724
rect 27648 44788 27738 44800
rect 27648 44724 27660 44788
rect 27724 44724 27738 44788
rect 27648 44710 27738 44724
rect 28200 44788 28290 44800
rect 28200 44724 28212 44788
rect 28276 44724 28290 44788
rect 28200 44710 28290 44724
rect 28752 44788 28842 44800
rect 28752 44724 28764 44788
rect 28828 44724 28842 44788
rect 28752 44710 28842 44724
rect 29304 44788 29394 44800
rect 29304 44724 29316 44788
rect 29380 44724 29394 44788
rect 29304 44710 29394 44724
rect 200 6655 600 44400
rect 1600 44300 2400 44400
rect 800 43300 1200 44152
rect 1600 43600 65400 44300
rect 4400 43300 5300 43400
rect 800 42800 4500 43300
rect 5200 42800 5300 43300
rect 199 6654 601 6655
rect 199 6254 200 6654
rect 600 6254 601 6654
rect 199 6253 601 6254
rect 200 1000 600 6253
rect 800 6134 1200 42800
rect 4400 42700 5300 42800
rect 5728 41840 6048 43600
rect 6300 43300 6800 43400
rect 6300 42800 6400 43300
rect 6700 42800 6800 43300
rect 6300 42700 6800 42800
rect 6388 42026 6708 42700
rect 13502 41740 13822 43600
rect 14074 43300 14574 43400
rect 14074 42800 14174 43300
rect 14474 42800 14574 43300
rect 14074 42700 14574 42800
rect 14162 42026 14482 42700
rect 21276 41640 21596 43600
rect 21848 43300 22348 43400
rect 21848 42800 21948 43300
rect 22248 42800 22348 43300
rect 21848 42700 22348 42800
rect 21936 42026 22256 42700
rect 29050 41540 29370 43600
rect 29622 43300 30122 43400
rect 29622 42800 29722 43300
rect 30022 42800 30122 43300
rect 29622 42700 30122 42800
rect 29710 42026 30030 42700
rect 36824 41540 37144 43600
rect 37396 43300 37896 43400
rect 37396 42800 37496 43300
rect 37796 42800 37896 43300
rect 37396 42700 37896 42800
rect 37484 42026 37804 42700
rect 44598 41540 44918 43600
rect 45170 43300 45670 43400
rect 45170 42800 45270 43300
rect 45570 42800 45670 43300
rect 45170 42700 45670 42800
rect 45258 42026 45578 42700
rect 52372 41540 52692 43600
rect 52944 43300 53444 43400
rect 52944 42800 53044 43300
rect 53344 42800 53444 43300
rect 52944 42700 53444 42800
rect 53032 42026 53352 42700
rect 60146 41540 60466 43600
rect 60718 43300 61218 43400
rect 60718 42800 60818 43300
rect 61118 42800 61218 43300
rect 60718 42700 61218 42800
rect 60806 42026 61126 42700
rect 1520 6653 25558 6654
rect 1520 6255 1521 6653
rect 1919 6255 25558 6653
rect 1520 6254 25558 6255
rect 800 5734 25558 6134
rect 800 1000 1200 5734
rect 5780 5089 6020 5120
rect 5780 4911 5811 5089
rect 5989 4911 6020 5089
rect 5780 4880 6020 4911
rect 5810 890 5990 4880
rect 21122 3299 24120 3300
rect 11432 3289 11752 3290
rect 11432 2971 11433 3289
rect 11751 2971 11752 3289
rect 21122 3009 21123 3299
rect 21413 3009 24120 3299
rect 21122 3008 24120 3009
rect 30785 3240 31063 3241
rect 11432 1916 11752 2971
rect 23884 2218 24064 3008
rect 30785 2964 30786 3240
rect 31062 2964 31063 3240
rect 23884 2038 26678 2218
rect 11432 1736 22814 1916
rect 11432 1666 11752 1736
rect 5810 710 18950 890
rect 3314 0 3494 200
rect 7178 0 7358 200
rect 11042 0 11222 200
rect 14906 0 15086 200
rect 18770 0 18950 710
rect 22634 0 22814 1736
rect 26498 0 26678 2038
rect 30785 1634 31063 2964
rect 30362 1454 31063 1634
rect 30362 0 30542 1454
rect 30785 1405 31063 1454
rect 65000 1000 65400 43600
rect 65600 43400 66000 44152
rect 65600 43300 66100 43400
rect 65600 42800 65700 43300
rect 66000 42800 66100 43300
rect 65600 42700 66100 42800
rect 65600 1000 66000 42700
use analog_control_wrapper  analog_control_wrapper_1
timestamp 1740731205
transform 1 0 2072 0 1 2042
box 514 496 62414 41000
use segdac  segdac_0
timestamp 1725599052
transform 1 0 27099 0 1 3114
box -1901 -360 4160 5600
use segdac  segdac_blue
timestamp 1725599052
transform 1 0 7779 0 1 3114
box -1901 -360 4160 5600
use segdac  segdac_green
timestamp 1725599052
transform 1 0 17439 0 1 3114
box -1901 -360 4160 5600
<< labels >>
flabel metal4 s 28766 44952 28826 45152 0 FreeSans 480 90 0 0 clk
port 0 nsew signal input
flabel metal4 s 29318 44952 29378 45152 0 FreeSans 480 90 0 0 ena
port 1 nsew signal input
flabel metal4 s 28214 44952 28274 45152 0 FreeSans 480 90 0 0 rst_n
port 2 nsew signal input
flabel metal4 s 30362 0 30542 200 0 FreeSans 960 0 0 0 ua[0]
port 3 nsew signal bidirectional
flabel metal4 s 26498 0 26678 200 0 FreeSans 960 0 0 0 ua[1]
port 4 nsew signal bidirectional
flabel metal4 s 22634 0 22814 200 0 FreeSans 960 0 0 0 ua[2]
port 5 nsew signal bidirectional
flabel metal4 s 18770 0 18950 200 0 FreeSans 960 0 0 0 ua[3]
port 6 nsew signal bidirectional
flabel metal4 s 14906 0 15086 200 0 FreeSans 960 0 0 0 ua[4]
port 7 nsew signal bidirectional
flabel metal4 s 11042 0 11222 200 0 FreeSans 960 0 0 0 ua[5]
port 8 nsew signal bidirectional
flabel metal4 s 7178 0 7358 200 0 FreeSans 960 0 0 0 ua[6]
port 9 nsew signal bidirectional
flabel metal4 s 3314 0 3494 200 0 FreeSans 960 0 0 0 ua[7]
port 10 nsew signal bidirectional
flabel metal4 s 27662 44952 27722 45152 0 FreeSans 480 90 0 0 ui_in[0]
port 11 nsew signal input
flabel metal4 s 27110 44952 27170 45152 0 FreeSans 480 90 0 0 ui_in[1]
port 12 nsew signal input
flabel metal4 s 26558 44952 26618 45152 0 FreeSans 480 90 0 0 ui_in[2]
port 13 nsew signal input
flabel metal4 s 26006 44952 26066 45152 0 FreeSans 480 90 0 0 ui_in[3]
port 14 nsew signal input
flabel metal4 s 25454 44952 25514 45152 0 FreeSans 480 90 0 0 ui_in[4]
port 15 nsew signal input
flabel metal4 s 24902 44952 24962 45152 0 FreeSans 480 90 0 0 ui_in[5]
port 16 nsew signal input
flabel metal4 s 24350 44952 24410 45152 0 FreeSans 480 90 0 0 ui_in[6]
port 17 nsew signal input
flabel metal4 s 23798 44952 23858 45152 0 FreeSans 480 90 0 0 ui_in[7]
port 18 nsew signal input
flabel metal4 s 23246 44952 23306 45152 0 FreeSans 480 90 0 0 uio_in[0]
port 19 nsew signal input
flabel metal4 s 22694 44952 22754 45152 0 FreeSans 480 90 0 0 uio_in[1]
port 20 nsew signal input
flabel metal4 s 22142 44952 22202 45152 0 FreeSans 480 90 0 0 uio_in[2]
port 21 nsew signal input
flabel metal4 s 21590 44952 21650 45152 0 FreeSans 480 90 0 0 uio_in[3]
port 22 nsew signal input
flabel metal4 s 21038 44952 21098 45152 0 FreeSans 480 90 0 0 uio_in[4]
port 23 nsew signal input
flabel metal4 s 20486 44952 20546 45152 0 FreeSans 480 90 0 0 uio_in[5]
port 24 nsew signal input
flabel metal4 s 19934 44952 19994 45152 0 FreeSans 480 90 0 0 uio_in[6]
port 25 nsew signal input
flabel metal4 s 19382 44952 19442 45152 0 FreeSans 480 90 0 0 uio_in[7]
port 26 nsew signal input
flabel metal4 s 9998 44952 10058 45152 0 FreeSans 480 90 0 0 uio_oe[0]
port 27 nsew signal output
flabel metal4 s 9446 44952 9506 45152 0 FreeSans 480 90 0 0 uio_oe[1]
port 28 nsew signal output
flabel metal4 s 8894 44952 8954 45152 0 FreeSans 480 90 0 0 uio_oe[2]
port 29 nsew signal output
flabel metal4 s 8342 44952 8402 45152 0 FreeSans 480 90 0 0 uio_oe[3]
port 30 nsew signal output
flabel metal4 s 7790 44952 7850 45152 0 FreeSans 480 90 0 0 uio_oe[4]
port 31 nsew signal output
flabel metal4 s 7238 44952 7298 45152 0 FreeSans 480 90 0 0 uio_oe[5]
port 32 nsew signal output
flabel metal4 s 6686 44952 6746 45152 0 FreeSans 480 90 0 0 uio_oe[6]
port 33 nsew signal output
flabel metal4 s 6134 44952 6194 45152 0 FreeSans 480 90 0 0 uio_oe[7]
port 34 nsew signal output
flabel metal4 s 14414 44952 14474 45152 0 FreeSans 480 90 0 0 uio_out[0]
port 35 nsew signal output
flabel metal4 s 13862 44952 13922 45152 0 FreeSans 480 90 0 0 uio_out[1]
port 36 nsew signal output
flabel metal4 s 13310 44952 13370 45152 0 FreeSans 480 90 0 0 uio_out[2]
port 37 nsew signal output
flabel metal4 s 12758 44952 12818 45152 0 FreeSans 480 90 0 0 uio_out[3]
port 38 nsew signal output
flabel metal4 s 12206 44952 12266 45152 0 FreeSans 480 90 0 0 uio_out[4]
port 39 nsew signal output
flabel metal4 s 11654 44952 11714 45152 0 FreeSans 480 90 0 0 uio_out[5]
port 40 nsew signal output
flabel metal4 s 11102 44952 11162 45152 0 FreeSans 480 90 0 0 uio_out[6]
port 41 nsew signal output
flabel metal4 s 10550 44952 10610 45152 0 FreeSans 480 90 0 0 uio_out[7]
port 42 nsew signal output
flabel metal4 s 18830 44952 18890 45152 0 FreeSans 480 90 0 0 uo_out[0]
port 43 nsew signal output
flabel metal4 s 18278 44952 18338 45152 0 FreeSans 480 90 0 0 uo_out[1]
port 44 nsew signal output
flabel metal4 s 17726 44952 17786 45152 0 FreeSans 480 90 0 0 uo_out[2]
port 45 nsew signal output
flabel metal4 s 17174 44952 17234 45152 0 FreeSans 480 90 0 0 uo_out[3]
port 46 nsew signal output
flabel metal4 s 16622 44952 16682 45152 0 FreeSans 480 90 0 0 uo_out[4]
port 47 nsew signal output
flabel metal4 s 16070 44952 16130 45152 0 FreeSans 480 90 0 0 uo_out[5]
port 48 nsew signal output
flabel metal4 s 15518 44952 15578 45152 0 FreeSans 480 90 0 0 uo_out[6]
port 49 nsew signal output
flabel metal4 s 14966 44952 15026 45152 0 FreeSans 480 90 0 0 uo_out[7]
port 50 nsew signal output
flabel metal4 200 1000 600 44152 1 FreeSans 400 0 0 0 VDPWR
port 51 nsew power bidirectional
flabel metal4 800 1000 1200 44152 1 FreeSans 400 0 0 0 VGND
port 52 nsew ground bidirectional
flabel metal4 65000 1000 65400 44152 1 FreeSans 400 0 0 0 VDPWR
port 51 nsew power bidirectional
flabel metal4 65600 1000 66000 44152 1 FreeSans 400 0 0 0 VGND
port 52 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 66976 45152
<< end >>
